library ieee;
use ieee.std_logic_1164.all;

entity ent is
    port (
         : in std_logic;
        rst : in std_logic;
        sig
    );
end ent;

architecture rtl of ent is

begin

end architecture;